

package axi4lite_pkg;

  `include "axi4lite_base.svh"
  `include "Axi4lite_Transaction.svh"
  // `include "axi4_monitor.svh"
  `include "axi4lite_master.svh"
  // `include "axi4_slave.svh"

endpackage