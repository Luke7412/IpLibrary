


interface UartIntf();

  logic rx;
  logic tx;
  string state;

endinterface