

package axi4s_pkg;

  `include "axi4s_base.svh"
  `include "axi4s_monitor.svh"
  `include "axi4s_master.svh"
  `include "axi4s_slave.svh"

endpackage