
--------------------------------------------------------------------------------
-- Info
--------------------------------------------------------------------------------
-- Hash (MD5): 0xf8e09f8403f237056f65015958b2728b
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- LIBRARIES
--------------------------------------------------------------------------------
library IEEE;
   use IEEE.STD_LOGIC_1164.ALL;


--------------------------------------------------------------------------------
-- PACKAGE HEADER
--------------------------------------------------------------------------------
package ModuleId is
   
   constant Id : std_logic_vector(127 downto 0) := X"f8e09f8403f237056f65015958b2728b";

end package;