

package types_pkg;

  typedef logic [ 7:0] u8;
  typedef logic [15:0] u16;
  typedef logic [31:0] u32;
  typedef logic [31:0] u64;

  typedef signed logic [ 7:0] i8;
  typedef signed logic [15:0] i16;
  typedef signed logic [31:0] i32;
  typedef signed logic [31:0] i64;

endpackage