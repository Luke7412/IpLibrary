//------------------------------------------------------------------------------
// Project Name: IpLibrary
//------------------------------------------------------------------------------
// Author      : Lukas Vinkx (lvin)
// Description : 
//------------------------------------------------------------------------------


`timescale 1ns/1ns;


package uart_pkg;

  `include "uart_base.svh";
  `include "uart_transmitter.svh";
  `include "uart_receiver.svh";

endpackage