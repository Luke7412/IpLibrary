
package coding_8b10b_pkg;


  typedef struct {
    string name;
    logic [7:0] code_8b;
    logic is_k;
    logic [9:0] code_10b_n;
    logic [9:0] code_10b_p;
    logic flip_rd;
  } t_entry;


  localparam t_entry entries [] = '{
  // {name: "Dx.y" , is_k: ?  code_8b:   HGF_EDCBA, code_10b_p:   jhgf_iedcba, code_10b_n:   jhgf_iedcba, flip_rd: ?} ,
    '{name: "D0.0" , is_k: 0, code_8b: 'b000_00000, code_10b_p: 'b0010_111001, code_10b_n: 'b1101_000110, flip_rd: 0},
    '{name: "D0.1" , is_k: 0, code_8b: 'b001_00000, code_10b_p: 'b1001_111001, code_10b_n: 'b1001_000110, flip_rd: 1},
    '{name: "D0.2" , is_k: 0, code_8b: 'b010_00000, code_10b_p: 'b1010_111001, code_10b_n: 'b1010_000110, flip_rd: 1},
    '{name: "D0.3" , is_k: 0, code_8b: 'b011_00000, code_10b_p: 'b1100_111001, code_10b_n: 'b0011_000110, flip_rd: 1},
    '{name: "D0.4" , is_k: 0, code_8b: 'b100_00000, code_10b_p: 'b0100_111001, code_10b_n: 'b1011_000110, flip_rd: 0},
    '{name: "D0.5" , is_k: 0, code_8b: 'b101_00000, code_10b_p: 'b0101_111001, code_10b_n: 'b0101_000110, flip_rd: 1},
    '{name: "D0.6" , is_k: 0, code_8b: 'b110_00000, code_10b_p: 'b0110_111001, code_10b_n: 'b0110_000110, flip_rd: 1},
    '{name: "D0.7" , is_k: 0, code_8b: 'b111_00000, code_10b_p: 'b1000_111001, code_10b_n: 'b0111_000110, flip_rd: 0},
    '{name: "D1.0" , is_k: 0, code_8b: 'b000_00001, code_10b_p: 'b0010_101110, code_10b_n: 'b1101_010001, flip_rd: 0},
    '{name: "D1.1" , is_k: 0, code_8b: 'b001_00001, code_10b_p: 'b1001_101110, code_10b_n: 'b1001_010001, flip_rd: 1},
    '{name: "D1.2" , is_k: 0, code_8b: 'b010_00001, code_10b_p: 'b1010_101110, code_10b_n: 'b1010_010001, flip_rd: 1},
    '{name: "D1.3" , is_k: 0, code_8b: 'b011_00001, code_10b_p: 'b1100_101110, code_10b_n: 'b0011_010001, flip_rd: 1},
    '{name: "D1.4" , is_k: 0, code_8b: 'b100_00001, code_10b_p: 'b0100_101110, code_10b_n: 'b1011_010001, flip_rd: 0},
    '{name: "D1.5" , is_k: 0, code_8b: 'b101_00001, code_10b_p: 'b0101_101110, code_10b_n: 'b0101_010001, flip_rd: 1},
    '{name: "D1.6" , is_k: 0, code_8b: 'b110_00001, code_10b_p: 'b0110_101110, code_10b_n: 'b0110_010001, flip_rd: 1},
    '{name: "D1.7" , is_k: 0, code_8b: 'b111_00001, code_10b_p: 'b1000_101110, code_10b_n: 'b0111_010001, flip_rd: 0},
    '{name: "D2.0" , is_k: 0, code_8b: 'b000_00010, code_10b_p: 'b0010_101101, code_10b_n: 'b1101_010010, flip_rd: 0},
    '{name: "D2.1" , is_k: 0, code_8b: 'b001_00010, code_10b_p: 'b1001_101101, code_10b_n: 'b1001_010010, flip_rd: 1},
    '{name: "D2.2" , is_k: 0, code_8b: 'b010_00010, code_10b_p: 'b1010_101101, code_10b_n: 'b1010_010010, flip_rd: 1},
    '{name: "D2.3" , is_k: 0, code_8b: 'b011_00010, code_10b_p: 'b1100_101101, code_10b_n: 'b0011_010010, flip_rd: 1},
    '{name: "D2.4" , is_k: 0, code_8b: 'b100_00010, code_10b_p: 'b0100_101101, code_10b_n: 'b1011_010010, flip_rd: 0},
    '{name: "D2.5" , is_k: 0, code_8b: 'b101_00010, code_10b_p: 'b0101_101101, code_10b_n: 'b0101_010010, flip_rd: 1},
    '{name: "D2.6" , is_k: 0, code_8b: 'b110_00010, code_10b_p: 'b0110_101101, code_10b_n: 'b0110_010010, flip_rd: 1},
    '{name: "D2.7" , is_k: 0, code_8b: 'b111_00010, code_10b_p: 'b1000_101101, code_10b_n: 'b0111_010010, flip_rd: 0},
    '{name: "D3.0" , is_k: 0, code_8b: 'b000_00011, code_10b_p: 'b1101_100011, code_10b_n: 'b0010_100011, flip_rd: 1},
    '{name: "D3.1" , is_k: 0, code_8b: 'b001_00011, code_10b_p: 'b1001_100011, code_10b_n: 'b1001_100011, flip_rd: 0},
    '{name: "D3.2" , is_k: 0, code_8b: 'b010_00011, code_10b_p: 'b1010_100011, code_10b_n: 'b1010_100011, flip_rd: 0},
    '{name: "D3.3" , is_k: 0, code_8b: 'b011_00011, code_10b_p: 'b0011_100011, code_10b_n: 'b1100_100011, flip_rd: 0},
    '{name: "D3.4" , is_k: 0, code_8b: 'b100_00011, code_10b_p: 'b1011_100011, code_10b_n: 'b0100_100011, flip_rd: 1},
    '{name: "D3.5" , is_k: 0, code_8b: 'b101_00011, code_10b_p: 'b0101_100011, code_10b_n: 'b0101_100011, flip_rd: 0},
    '{name: "D3.6" , is_k: 0, code_8b: 'b110_00011, code_10b_p: 'b0110_100011, code_10b_n: 'b0110_100011, flip_rd: 0},
    '{name: "D3.7" , is_k: 0, code_8b: 'b111_00011, code_10b_p: 'b0111_100011, code_10b_n: 'b1000_100011, flip_rd: 1},
    '{name: "D4.0" , is_k: 0, code_8b: 'b000_00100, code_10b_p: 'b0010_101011, code_10b_n: 'b1101_010100, flip_rd: 0},
    '{name: "D4.1" , is_k: 0, code_8b: 'b001_00100, code_10b_p: 'b1001_101011, code_10b_n: 'b1001_010100, flip_rd: 1},
    '{name: "D4.2" , is_k: 0, code_8b: 'b010_00100, code_10b_p: 'b1010_101011, code_10b_n: 'b1010_010100, flip_rd: 1},
    '{name: "D4.3" , is_k: 0, code_8b: 'b011_00100, code_10b_p: 'b1100_101011, code_10b_n: 'b0011_010100, flip_rd: 1},
    '{name: "D4.4" , is_k: 0, code_8b: 'b100_00100, code_10b_p: 'b0100_101011, code_10b_n: 'b1011_010100, flip_rd: 0},
    '{name: "D4.5" , is_k: 0, code_8b: 'b101_00100, code_10b_p: 'b0101_101011, code_10b_n: 'b0101_010100, flip_rd: 1},
    '{name: "D4.6" , is_k: 0, code_8b: 'b110_00100, code_10b_p: 'b0110_101011, code_10b_n: 'b0110_010100, flip_rd: 1},
    '{name: "D4.7" , is_k: 0, code_8b: 'b111_00100, code_10b_p: 'b1000_101011, code_10b_n: 'b0111_010100, flip_rd: 0},
    '{name: "D5.0" , is_k: 0, code_8b: 'b000_00101, code_10b_p: 'b1101_100101, code_10b_n: 'b0010_100101, flip_rd: 1},
    '{name: "D5.1" , is_k: 0, code_8b: 'b001_00101, code_10b_p: 'b1001_100101, code_10b_n: 'b1001_100101, flip_rd: 0},
    '{name: "D5.2" , is_k: 0, code_8b: 'b010_00101, code_10b_p: 'b1010_100101, code_10b_n: 'b1010_100101, flip_rd: 0},
    '{name: "D5.3" , is_k: 0, code_8b: 'b011_00101, code_10b_p: 'b0011_100101, code_10b_n: 'b1100_100101, flip_rd: 0},
    '{name: "D5.4" , is_k: 0, code_8b: 'b100_00101, code_10b_p: 'b1011_100101, code_10b_n: 'b0100_100101, flip_rd: 1},
    '{name: "D5.5" , is_k: 0, code_8b: 'b101_00101, code_10b_p: 'b0101_100101, code_10b_n: 'b0101_100101, flip_rd: 0},
    '{name: "D5.6" , is_k: 0, code_8b: 'b110_00101, code_10b_p: 'b0110_100101, code_10b_n: 'b0110_100101, flip_rd: 0},
    '{name: "D5.7" , is_k: 0, code_8b: 'b111_00101, code_10b_p: 'b0111_100101, code_10b_n: 'b1000_100101, flip_rd: 1},
    '{name: "D6.0" , is_k: 0, code_8b: 'b000_00110, code_10b_p: 'b1101_100110, code_10b_n: 'b0010_100110, flip_rd: 1},
    '{name: "D6.1" , is_k: 0, code_8b: 'b001_00110, code_10b_p: 'b1001_100110, code_10b_n: 'b1001_100110, flip_rd: 0},
    '{name: "D6.2" , is_k: 0, code_8b: 'b010_00110, code_10b_p: 'b1010_100110, code_10b_n: 'b1010_100110, flip_rd: 0},
    '{name: "D6.3" , is_k: 0, code_8b: 'b011_00110, code_10b_p: 'b0011_100110, code_10b_n: 'b1100_100110, flip_rd: 0},
    '{name: "D6.4" , is_k: 0, code_8b: 'b100_00110, code_10b_p: 'b1011_100110, code_10b_n: 'b0100_100110, flip_rd: 1},
    '{name: "D6.5" , is_k: 0, code_8b: 'b101_00110, code_10b_p: 'b0101_100110, code_10b_n: 'b0101_100110, flip_rd: 0},
    '{name: "D6.6" , is_k: 0, code_8b: 'b110_00110, code_10b_p: 'b0110_100110, code_10b_n: 'b0110_100110, flip_rd: 0},
    '{name: "D6.7" , is_k: 0, code_8b: 'b111_00110, code_10b_p: 'b0111_100110, code_10b_n: 'b1000_100110, flip_rd: 1},
    '{name: "D7.0" , is_k: 0, code_8b: 'b000_00111, code_10b_p: 'b1101_000111, code_10b_n: 'b0010_111000, flip_rd: 1},
    '{name: "D7.1" , is_k: 0, code_8b: 'b001_00111, code_10b_p: 'b1001_000111, code_10b_n: 'b1001_111000, flip_rd: 0},
    '{name: "D7.2" , is_k: 0, code_8b: 'b010_00111, code_10b_p: 'b1010_000111, code_10b_n: 'b1010_111000, flip_rd: 0},
    '{name: "D7.3" , is_k: 0, code_8b: 'b011_00111, code_10b_p: 'b0011_000111, code_10b_n: 'b1100_111000, flip_rd: 0},
    '{name: "D7.4" , is_k: 0, code_8b: 'b100_00111, code_10b_p: 'b1011_000111, code_10b_n: 'b0100_111000, flip_rd: 1},
    '{name: "D7.5" , is_k: 0, code_8b: 'b101_00111, code_10b_p: 'b0101_000111, code_10b_n: 'b0101_111000, flip_rd: 0},
    '{name: "D7.6" , is_k: 0, code_8b: 'b110_00111, code_10b_p: 'b0110_000111, code_10b_n: 'b0110_111000, flip_rd: 0},
    '{name: "D7.7" , is_k: 0, code_8b: 'b111_00111, code_10b_p: 'b0111_000111, code_10b_n: 'b1000_111000, flip_rd: 1},
    '{name: "D8.0" , is_k: 0, code_8b: 'b000_01000, code_10b_p: 'b0010_100111, code_10b_n: 'b1101_011000, flip_rd: 0},
    '{name: "D8.1" , is_k: 0, code_8b: 'b001_01000, code_10b_p: 'b1001_100111, code_10b_n: 'b1001_011000, flip_rd: 1},
    '{name: "D8.2" , is_k: 0, code_8b: 'b010_01000, code_10b_p: 'b1010_100111, code_10b_n: 'b1010_011000, flip_rd: 1},
    '{name: "D8.3" , is_k: 0, code_8b: 'b011_01000, code_10b_p: 'b1100_100111, code_10b_n: 'b0011_011000, flip_rd: 1},
    '{name: "D8.4" , is_k: 0, code_8b: 'b100_01000, code_10b_p: 'b0100_100111, code_10b_n: 'b1011_011000, flip_rd: 0},
    '{name: "D8.5" , is_k: 0, code_8b: 'b101_01000, code_10b_p: 'b0101_100111, code_10b_n: 'b0101_011000, flip_rd: 1},
    '{name: "D8.6" , is_k: 0, code_8b: 'b110_01000, code_10b_p: 'b0110_100111, code_10b_n: 'b0110_011000, flip_rd: 1},
    '{name: "D8.7" , is_k: 0, code_8b: 'b111_01000, code_10b_p: 'b1000_100111, code_10b_n: 'b0111_011000, flip_rd: 0},
    '{name: "D9.0" , is_k: 0, code_8b: 'b000_01001, code_10b_p: 'b1101_101001, code_10b_n: 'b0010_101001, flip_rd: 1},
    '{name: "D9.1" , is_k: 0, code_8b: 'b001_01001, code_10b_p: 'b1001_101001, code_10b_n: 'b1001_101001, flip_rd: 0},
    '{name: "D9.2" , is_k: 0, code_8b: 'b010_01001, code_10b_p: 'b1010_101001, code_10b_n: 'b1010_101001, flip_rd: 0},
    '{name: "D9.3" , is_k: 0, code_8b: 'b011_01001, code_10b_p: 'b0011_101001, code_10b_n: 'b1100_101001, flip_rd: 0},
    '{name: "D9.4" , is_k: 0, code_8b: 'b100_01001, code_10b_p: 'b1011_101001, code_10b_n: 'b0100_101001, flip_rd: 1},
    '{name: "D9.5" , is_k: 0, code_8b: 'b101_01001, code_10b_p: 'b0101_101001, code_10b_n: 'b0101_101001, flip_rd: 0},
    '{name: "D9.6" , is_k: 0, code_8b: 'b110_01001, code_10b_p: 'b0110_101001, code_10b_n: 'b0110_101001, flip_rd: 0},
    '{name: "D9.7" , is_k: 0, code_8b: 'b111_01001, code_10b_p: 'b0111_101001, code_10b_n: 'b1000_101001, flip_rd: 1},
    '{name: "D10.0", is_k: 0, code_8b: 'b000_01010, code_10b_p: 'b1101_101010, code_10b_n: 'b0010_101010, flip_rd: 1},
    '{name: "D10.1", is_k: 0, code_8b: 'b001_01010, code_10b_p: 'b1001_101010, code_10b_n: 'b1001_101010, flip_rd: 0},
    '{name: "D10.2", is_k: 0, code_8b: 'b010_01010, code_10b_p: 'b1010_101010, code_10b_n: 'b1010_101010, flip_rd: 0},
    '{name: "D10.3", is_k: 0, code_8b: 'b011_01010, code_10b_p: 'b0011_101010, code_10b_n: 'b1100_101010, flip_rd: 0},
    '{name: "D10.4", is_k: 0, code_8b: 'b100_01010, code_10b_p: 'b1011_101010, code_10b_n: 'b0100_101010, flip_rd: 1},
    '{name: "D10.5", is_k: 0, code_8b: 'b101_01010, code_10b_p: 'b0101_101010, code_10b_n: 'b0101_101010, flip_rd: 0},
    '{name: "D10.6", is_k: 0, code_8b: 'b110_01010, code_10b_p: 'b0110_101010, code_10b_n: 'b0110_101010, flip_rd: 0},
    '{name: "D10.7", is_k: 0, code_8b: 'b111_01010, code_10b_p: 'b0111_101010, code_10b_n: 'b1000_101010, flip_rd: 1},
    '{name: "D11.0", is_k: 0, code_8b: 'b000_01011, code_10b_p: 'b1101_001011, code_10b_n: 'b0010_001011, flip_rd: 1},
    '{name: "D11.1", is_k: 0, code_8b: 'b001_01011, code_10b_p: 'b1001_001011, code_10b_n: 'b1001_001011, flip_rd: 0},
    '{name: "D11.2", is_k: 0, code_8b: 'b010_01011, code_10b_p: 'b1010_001011, code_10b_n: 'b1010_001011, flip_rd: 0},
    '{name: "D11.3", is_k: 0, code_8b: 'b011_01011, code_10b_p: 'b0011_001011, code_10b_n: 'b1100_001011, flip_rd: 0},
    '{name: "D11.4", is_k: 0, code_8b: 'b100_01011, code_10b_p: 'b1011_001011, code_10b_n: 'b0100_001011, flip_rd: 1},
    '{name: "D11.5", is_k: 0, code_8b: 'b101_01011, code_10b_p: 'b0101_001011, code_10b_n: 'b0101_001011, flip_rd: 0},
    '{name: "D11.6", is_k: 0, code_8b: 'b110_01011, code_10b_p: 'b0110_001011, code_10b_n: 'b0110_001011, flip_rd: 0},
    '{name: "D11.7", is_k: 0, code_8b: 'b111_01011, code_10b_p: 'b0111_001011, code_10b_n: 'b0001_001011, flip_rd: 1},
    '{name: "D12.0", is_k: 0, code_8b: 'b000_01100, code_10b_p: 'b1101_101100, code_10b_n: 'b0010_101100, flip_rd: 1},
    '{name: "D12.1", is_k: 0, code_8b: 'b001_01100, code_10b_p: 'b1001_101100, code_10b_n: 'b1001_101100, flip_rd: 0},
    '{name: "D12.2", is_k: 0, code_8b: 'b010_01100, code_10b_p: 'b1010_101100, code_10b_n: 'b1010_101100, flip_rd: 0},
    '{name: "D12.3", is_k: 0, code_8b: 'b011_01100, code_10b_p: 'b0011_101100, code_10b_n: 'b1100_101100, flip_rd: 0},
    '{name: "D12.4", is_k: 0, code_8b: 'b100_01100, code_10b_p: 'b1011_101100, code_10b_n: 'b0100_101100, flip_rd: 1},
    '{name: "D12.5", is_k: 0, code_8b: 'b101_01100, code_10b_p: 'b0101_101100, code_10b_n: 'b0101_101100, flip_rd: 0},
    '{name: "D12.6", is_k: 0, code_8b: 'b110_01100, code_10b_p: 'b0110_101100, code_10b_n: 'b0110_101100, flip_rd: 0},
    '{name: "D12.7", is_k: 0, code_8b: 'b111_01100, code_10b_p: 'b0111_101100, code_10b_n: 'b1000_101100, flip_rd: 1},
    '{name: "D13.0", is_k: 0, code_8b: 'b000_01101, code_10b_p: 'b1101_001101, code_10b_n: 'b0010_001101, flip_rd: 1},
    '{name: "D13.1", is_k: 0, code_8b: 'b001_01101, code_10b_p: 'b1001_001101, code_10b_n: 'b1001_001101, flip_rd: 0},
    '{name: "D13.2", is_k: 0, code_8b: 'b010_01101, code_10b_p: 'b1010_001101, code_10b_n: 'b1010_001101, flip_rd: 0},
    '{name: "D13.3", is_k: 0, code_8b: 'b011_01101, code_10b_p: 'b0011_001101, code_10b_n: 'b1100_001101, flip_rd: 0},
    '{name: "D13.4", is_k: 0, code_8b: 'b100_01101, code_10b_p: 'b1011_001101, code_10b_n: 'b0100_001101, flip_rd: 1},
    '{name: "D13.5", is_k: 0, code_8b: 'b101_01101, code_10b_p: 'b0101_001101, code_10b_n: 'b0101_001101, flip_rd: 0},
    '{name: "D13.6", is_k: 0, code_8b: 'b110_01101, code_10b_p: 'b0110_001101, code_10b_n: 'b0110_001101, flip_rd: 0},
    '{name: "D13.7", is_k: 0, code_8b: 'b111_01101, code_10b_p: 'b0111_001101, code_10b_n: 'b0001_001101, flip_rd: 1},
    '{name: "D14.0", is_k: 0, code_8b: 'b000_01110, code_10b_p: 'b1101_001110, code_10b_n: 'b0010_001110, flip_rd: 1},
    '{name: "D14.1", is_k: 0, code_8b: 'b001_01110, code_10b_p: 'b1001_001110, code_10b_n: 'b1001_001110, flip_rd: 0},
    '{name: "D14.2", is_k: 0, code_8b: 'b010_01110, code_10b_p: 'b1010_001110, code_10b_n: 'b1010_001110, flip_rd: 0},
    '{name: "D14.3", is_k: 0, code_8b: 'b011_01110, code_10b_p: 'b0011_001110, code_10b_n: 'b1100_001110, flip_rd: 0},
    '{name: "D14.4", is_k: 0, code_8b: 'b100_01110, code_10b_p: 'b1011_001110, code_10b_n: 'b0100_001110, flip_rd: 1},
    '{name: "D14.5", is_k: 0, code_8b: 'b101_01110, code_10b_p: 'b0101_001110, code_10b_n: 'b0101_001110, flip_rd: 0},
    '{name: "D14.6", is_k: 0, code_8b: 'b110_01110, code_10b_p: 'b0110_001110, code_10b_n: 'b0110_001110, flip_rd: 0},
    '{name: "D14.7", is_k: 0, code_8b: 'b111_01110, code_10b_p: 'b0111_001110, code_10b_n: 'b0001_001110, flip_rd: 1},
    '{name: "D15.0", is_k: 0, code_8b: 'b000_01111, code_10b_p: 'b0010_111010, code_10b_n: 'b1101_000101, flip_rd: 0},
    '{name: "D15.1", is_k: 0, code_8b: 'b001_01111, code_10b_p: 'b1001_111010, code_10b_n: 'b1001_000101, flip_rd: 1},
    '{name: "D15.2", is_k: 0, code_8b: 'b010_01111, code_10b_p: 'b1010_111010, code_10b_n: 'b1010_000101, flip_rd: 1},
    '{name: "D15.3", is_k: 0, code_8b: 'b011_01111, code_10b_p: 'b1100_111010, code_10b_n: 'b0011_000101, flip_rd: 1},
    '{name: "D15.4", is_k: 0, code_8b: 'b100_01111, code_10b_p: 'b0100_111010, code_10b_n: 'b1011_000101, flip_rd: 0},
    '{name: "D15.5", is_k: 0, code_8b: 'b101_01111, code_10b_p: 'b0101_111010, code_10b_n: 'b0101_000101, flip_rd: 1},
    '{name: "D15.6", is_k: 0, code_8b: 'b110_01111, code_10b_p: 'b0110_111010, code_10b_n: 'b0110_000101, flip_rd: 1},
    '{name: "D15.7", is_k: 0, code_8b: 'b111_01111, code_10b_p: 'b1000_111010, code_10b_n: 'b0111_000101, flip_rd: 0},
    '{name: "D16.0", is_k: 0, code_8b: 'b000_10000, code_10b_p: 'b0010_110110, code_10b_n: 'b1101_001001, flip_rd: 0},
    '{name: "D16.1", is_k: 0, code_8b: 'b001_10000, code_10b_p: 'b1001_110110, code_10b_n: 'b1001_001001, flip_rd: 1},
    '{name: "D16.2", is_k: 0, code_8b: 'b010_10000, code_10b_p: 'b1010_110110, code_10b_n: 'b1010_001001, flip_rd: 1},
    '{name: "D16.3", is_k: 0, code_8b: 'b011_10000, code_10b_p: 'b1100_110110, code_10b_n: 'b0011_001001, flip_rd: 1},
    '{name: "D16.4", is_k: 0, code_8b: 'b100_10000, code_10b_p: 'b0100_110110, code_10b_n: 'b1011_001001, flip_rd: 0},
    '{name: "D16.5", is_k: 0, code_8b: 'b101_10000, code_10b_p: 'b0101_110110, code_10b_n: 'b0101_001001, flip_rd: 1},
    '{name: "D16.6", is_k: 0, code_8b: 'b110_10000, code_10b_p: 'b0110_110110, code_10b_n: 'b0110_001001, flip_rd: 1},
    '{name: "D16.7", is_k: 0, code_8b: 'b111_10000, code_10b_p: 'b1000_110110, code_10b_n: 'b0111_001001, flip_rd: 0},
    '{name: "D17.0", is_k: 0, code_8b: 'b000_10001, code_10b_p: 'b1101_110001, code_10b_n: 'b0010_110001, flip_rd: 1},
    '{name: "D17.1", is_k: 0, code_8b: 'b001_10001, code_10b_p: 'b1001_110001, code_10b_n: 'b1001_110001, flip_rd: 0},
    '{name: "D17.2", is_k: 0, code_8b: 'b010_10001, code_10b_p: 'b1010_110001, code_10b_n: 'b1010_110001, flip_rd: 0},
    '{name: "D17.3", is_k: 0, code_8b: 'b011_10001, code_10b_p: 'b0011_110001, code_10b_n: 'b1100_110001, flip_rd: 0},
    '{name: "D17.4", is_k: 0, code_8b: 'b100_10001, code_10b_p: 'b1011_110001, code_10b_n: 'b0100_110001, flip_rd: 1},
    '{name: "D17.5", is_k: 0, code_8b: 'b101_10001, code_10b_p: 'b0101_110001, code_10b_n: 'b0101_110001, flip_rd: 0},
    '{name: "D17.6", is_k: 0, code_8b: 'b110_10001, code_10b_p: 'b0110_110001, code_10b_n: 'b0110_110001, flip_rd: 0},
    '{name: "D17.7", is_k: 0, code_8b: 'b111_10001, code_10b_p: 'b1110_110001, code_10b_n: 'b1000_110001, flip_rd: 1},
    '{name: "D18.0", is_k: 0, code_8b: 'b000_10010, code_10b_p: 'b1101_110010, code_10b_n: 'b0010_110010, flip_rd: 1},
    '{name: "D18.1", is_k: 0, code_8b: 'b001_10010, code_10b_p: 'b1001_110010, code_10b_n: 'b1001_110010, flip_rd: 0},
    '{name: "D18.2", is_k: 0, code_8b: 'b010_10010, code_10b_p: 'b1010_110010, code_10b_n: 'b1010_110010, flip_rd: 0},
    '{name: "D18.3", is_k: 0, code_8b: 'b011_10010, code_10b_p: 'b0011_110010, code_10b_n: 'b1100_110010, flip_rd: 0},
    '{name: "D18.4", is_k: 0, code_8b: 'b100_10010, code_10b_p: 'b1011_110010, code_10b_n: 'b0100_110010, flip_rd: 1},
    '{name: "D18.5", is_k: 0, code_8b: 'b101_10010, code_10b_p: 'b0101_110010, code_10b_n: 'b0101_110010, flip_rd: 0},
    '{name: "D18.6", is_k: 0, code_8b: 'b110_10010, code_10b_p: 'b0110_110010, code_10b_n: 'b0110_110010, flip_rd: 0},
    '{name: "D18.7", is_k: 0, code_8b: 'b111_10010, code_10b_p: 'b1110_110010, code_10b_n: 'b1000_110010, flip_rd: 1},
    '{name: "D19.0", is_k: 0, code_8b: 'b000_10011, code_10b_p: 'b1101_010011, code_10b_n: 'b0010_010011, flip_rd: 1},
    '{name: "D19.1", is_k: 0, code_8b: 'b001_10011, code_10b_p: 'b1001_010011, code_10b_n: 'b1001_010011, flip_rd: 0},
    '{name: "D19.2", is_k: 0, code_8b: 'b010_10011, code_10b_p: 'b1010_010011, code_10b_n: 'b1010_010011, flip_rd: 0},
    '{name: "D19.3", is_k: 0, code_8b: 'b011_10011, code_10b_p: 'b0011_010011, code_10b_n: 'b1100_010011, flip_rd: 0},
    '{name: "D19.4", is_k: 0, code_8b: 'b100_10011, code_10b_p: 'b1011_010011, code_10b_n: 'b0100_010011, flip_rd: 1},
    '{name: "D19.5", is_k: 0, code_8b: 'b101_10011, code_10b_p: 'b0101_010011, code_10b_n: 'b0101_010011, flip_rd: 0},
    '{name: "D19.6", is_k: 0, code_8b: 'b110_10011, code_10b_p: 'b0110_010011, code_10b_n: 'b0110_010011, flip_rd: 0},
    '{name: "D19.7", is_k: 0, code_8b: 'b111_10011, code_10b_p: 'b0111_010011, code_10b_n: 'b1000_010011, flip_rd: 1},
    '{name: "D20.0", is_k: 0, code_8b: 'b000_10100, code_10b_p: 'b1101_110100, code_10b_n: 'b0010_110100, flip_rd: 1},
    '{name: "D20.1", is_k: 0, code_8b: 'b001_10100, code_10b_p: 'b1001_110100, code_10b_n: 'b1001_110100, flip_rd: 0},
    '{name: "D20.2", is_k: 0, code_8b: 'b010_10100, code_10b_p: 'b1010_110100, code_10b_n: 'b1010_110100, flip_rd: 0},
    '{name: "D20.3", is_k: 0, code_8b: 'b011_10100, code_10b_p: 'b0011_110100, code_10b_n: 'b1100_110100, flip_rd: 0},
    '{name: "D20.4", is_k: 0, code_8b: 'b100_10100, code_10b_p: 'b1011_110100, code_10b_n: 'b0100_110100, flip_rd: 1},
    '{name: "D20.5", is_k: 0, code_8b: 'b101_10100, code_10b_p: 'b0101_110100, code_10b_n: 'b0101_110100, flip_rd: 0},
    '{name: "D20.6", is_k: 0, code_8b: 'b110_10100, code_10b_p: 'b0110_110100, code_10b_n: 'b0110_110100, flip_rd: 0},
    '{name: "D20.7", is_k: 0, code_8b: 'b111_10100, code_10b_p: 'b1110_110100, code_10b_n: 'b1000_110100, flip_rd: 1},
    '{name: "D21.0", is_k: 0, code_8b: 'b000_10101, code_10b_p: 'b1101_010101, code_10b_n: 'b0010_010101, flip_rd: 1},
    '{name: "D21.1", is_k: 0, code_8b: 'b001_10101, code_10b_p: 'b1001_010101, code_10b_n: 'b1001_010101, flip_rd: 0},
    '{name: "D21.2", is_k: 0, code_8b: 'b010_10101, code_10b_p: 'b1010_010101, code_10b_n: 'b1010_010101, flip_rd: 0},
    '{name: "D21.3", is_k: 0, code_8b: 'b011_10101, code_10b_p: 'b0011_010101, code_10b_n: 'b1100_010101, flip_rd: 0},
    '{name: "D21.4", is_k: 0, code_8b: 'b100_10101, code_10b_p: 'b1011_010101, code_10b_n: 'b0100_010101, flip_rd: 1},
    '{name: "D21.5", is_k: 0, code_8b: 'b101_10101, code_10b_p: 'b0101_010101, code_10b_n: 'b0101_010101, flip_rd: 0},
    '{name: "D21.6", is_k: 0, code_8b: 'b110_10101, code_10b_p: 'b0110_010101, code_10b_n: 'b0110_010101, flip_rd: 0},
    '{name: "D21.7", is_k: 0, code_8b: 'b111_10101, code_10b_p: 'b0111_010101, code_10b_n: 'b1000_010101, flip_rd: 1},
    '{name: "D22.0", is_k: 0, code_8b: 'b000_10110, code_10b_p: 'b1101_010110, code_10b_n: 'b0010_010110, flip_rd: 1},
    '{name: "D22.1", is_k: 0, code_8b: 'b001_10110, code_10b_p: 'b1001_010110, code_10b_n: 'b1001_010110, flip_rd: 0},
    '{name: "D22.2", is_k: 0, code_8b: 'b010_10110, code_10b_p: 'b1010_010110, code_10b_n: 'b1010_010110, flip_rd: 0},
    '{name: "D22.3", is_k: 0, code_8b: 'b011_10110, code_10b_p: 'b0011_010110, code_10b_n: 'b1100_010110, flip_rd: 0},
    '{name: "D22.4", is_k: 0, code_8b: 'b100_10110, code_10b_p: 'b1011_010110, code_10b_n: 'b0100_010110, flip_rd: 1},
    '{name: "D22.5", is_k: 0, code_8b: 'b101_10110, code_10b_p: 'b0101_010110, code_10b_n: 'b0101_010110, flip_rd: 0},
    '{name: "D22.6", is_k: 0, code_8b: 'b110_10110, code_10b_p: 'b0110_010110, code_10b_n: 'b0110_010110, flip_rd: 0},
    '{name: "D22.7", is_k: 0, code_8b: 'b111_10110, code_10b_p: 'b0111_010110, code_10b_n: 'b1000_010110, flip_rd: 1},
    '{name: "D23.0", is_k: 0, code_8b: 'b000_10111, code_10b_p: 'b0010_010111, code_10b_n: 'b1101_101000, flip_rd: 0},
    '{name: "D23.1", is_k: 0, code_8b: 'b001_10111, code_10b_p: 'b1001_010111, code_10b_n: 'b1001_101000, flip_rd: 1},
    '{name: "D23.2", is_k: 0, code_8b: 'b010_10111, code_10b_p: 'b1010_010111, code_10b_n: 'b1010_101000, flip_rd: 1},
    '{name: "D23.3", is_k: 0, code_8b: 'b011_10111, code_10b_p: 'b1100_010111, code_10b_n: 'b0011_101000, flip_rd: 1},
    '{name: "D23.4", is_k: 0, code_8b: 'b100_10111, code_10b_p: 'b0100_010111, code_10b_n: 'b1011_101000, flip_rd: 0},
    '{name: "D23.5", is_k: 0, code_8b: 'b101_10111, code_10b_p: 'b0101_010111, code_10b_n: 'b0101_101000, flip_rd: 1},
    '{name: "D23.6", is_k: 0, code_8b: 'b110_10111, code_10b_p: 'b0110_010111, code_10b_n: 'b0110_101000, flip_rd: 1},
    '{name: "D23.7", is_k: 0, code_8b: 'b111_10111, code_10b_p: 'b1000_010111, code_10b_n: 'b0111_101000, flip_rd: 0},
    '{name: "D24.0", is_k: 0, code_8b: 'b000_11000, code_10b_p: 'b0010_110011, code_10b_n: 'b1101_001100, flip_rd: 0},
    '{name: "D24.1", is_k: 0, code_8b: 'b001_11000, code_10b_p: 'b1001_110011, code_10b_n: 'b1001_001100, flip_rd: 1},
    '{name: "D24.2", is_k: 0, code_8b: 'b010_11000, code_10b_p: 'b1010_110011, code_10b_n: 'b1010_001100, flip_rd: 1},
    '{name: "D24.3", is_k: 0, code_8b: 'b011_11000, code_10b_p: 'b1100_110011, code_10b_n: 'b0011_001100, flip_rd: 1},
    '{name: "D24.4", is_k: 0, code_8b: 'b100_11000, code_10b_p: 'b0100_110011, code_10b_n: 'b1011_001100, flip_rd: 0},
    '{name: "D24.5", is_k: 0, code_8b: 'b101_11000, code_10b_p: 'b0101_110011, code_10b_n: 'b0101_001100, flip_rd: 1},
    '{name: "D24.6", is_k: 0, code_8b: 'b110_11000, code_10b_p: 'b0110_110011, code_10b_n: 'b0110_001100, flip_rd: 1},
    '{name: "D24.7", is_k: 0, code_8b: 'b111_11000, code_10b_p: 'b1000_110011, code_10b_n: 'b0111_001100, flip_rd: 0},
    '{name: "D25.0", is_k: 0, code_8b: 'b000_11001, code_10b_p: 'b1101_011001, code_10b_n: 'b0010_011001, flip_rd: 1},
    '{name: "D25.1", is_k: 0, code_8b: 'b001_11001, code_10b_p: 'b1001_011001, code_10b_n: 'b1001_011001, flip_rd: 0},
    '{name: "D25.2", is_k: 0, code_8b: 'b010_11001, code_10b_p: 'b1010_011001, code_10b_n: 'b1010_011001, flip_rd: 0},
    '{name: "D25.3", is_k: 0, code_8b: 'b011_11001, code_10b_p: 'b0011_011001, code_10b_n: 'b1100_011001, flip_rd: 0},
    '{name: "D25.4", is_k: 0, code_8b: 'b100_11001, code_10b_p: 'b1011_011001, code_10b_n: 'b0100_011001, flip_rd: 1},
    '{name: "D25.5", is_k: 0, code_8b: 'b101_11001, code_10b_p: 'b0101_011001, code_10b_n: 'b0101_011001, flip_rd: 0},
    '{name: "D25.6", is_k: 0, code_8b: 'b110_11001, code_10b_p: 'b0110_011001, code_10b_n: 'b0110_011001, flip_rd: 0},
    '{name: "D25.7", is_k: 0, code_8b: 'b111_11001, code_10b_p: 'b0111_011001, code_10b_n: 'b1000_011001, flip_rd: 1},
    '{name: "D26.0", is_k: 0, code_8b: 'b000_11010, code_10b_p: 'b1101_011010, code_10b_n: 'b0010_011010, flip_rd: 1},
    '{name: "D26.1", is_k: 0, code_8b: 'b001_11010, code_10b_p: 'b1001_011010, code_10b_n: 'b1001_011010, flip_rd: 0},
    '{name: "D26.2", is_k: 0, code_8b: 'b010_11010, code_10b_p: 'b1010_011010, code_10b_n: 'b1010_011010, flip_rd: 0},
    '{name: "D26.3", is_k: 0, code_8b: 'b011_11010, code_10b_p: 'b0011_011010, code_10b_n: 'b1100_011010, flip_rd: 0},
    '{name: "D26.4", is_k: 0, code_8b: 'b100_11010, code_10b_p: 'b1011_011010, code_10b_n: 'b0100_011010, flip_rd: 1},
    '{name: "D26.5", is_k: 0, code_8b: 'b101_11010, code_10b_p: 'b0101_011010, code_10b_n: 'b0101_011010, flip_rd: 0},
    '{name: "D26.6", is_k: 0, code_8b: 'b110_11010, code_10b_p: 'b0110_011010, code_10b_n: 'b0110_011010, flip_rd: 0},
    '{name: "D26.7", is_k: 0, code_8b: 'b111_11010, code_10b_p: 'b0111_011010, code_10b_n: 'b1000_011010, flip_rd: 1},
    '{name: "D27.0", is_k: 0, code_8b: 'b000_11011, code_10b_p: 'b0010_011011, code_10b_n: 'b1101_100100, flip_rd: 0},
    '{name: "D27.1", is_k: 0, code_8b: 'b001_11011, code_10b_p: 'b1001_011011, code_10b_n: 'b1001_100100, flip_rd: 1},
    '{name: "D27.2", is_k: 0, code_8b: 'b010_11011, code_10b_p: 'b1010_011011, code_10b_n: 'b1010_100100, flip_rd: 1},
    '{name: "D27.3", is_k: 0, code_8b: 'b011_11011, code_10b_p: 'b1100_011011, code_10b_n: 'b0011_100100, flip_rd: 1},
    '{name: "D27.4", is_k: 0, code_8b: 'b100_11011, code_10b_p: 'b0100_011011, code_10b_n: 'b1011_100100, flip_rd: 0},
    '{name: "D27.5", is_k: 0, code_8b: 'b101_11011, code_10b_p: 'b0101_011011, code_10b_n: 'b0101_100100, flip_rd: 1},
    '{name: "D27.6", is_k: 0, code_8b: 'b110_11011, code_10b_p: 'b0110_011011, code_10b_n: 'b0110_100100, flip_rd: 1},
    '{name: "D27.7", is_k: 0, code_8b: 'b111_11011, code_10b_p: 'b1000_011011, code_10b_n: 'b0111_100100, flip_rd: 0},
    '{name: "D28.0", is_k: 0, code_8b: 'b000_11100, code_10b_p: 'b1101_011100, code_10b_n: 'b0010_011100, flip_rd: 1},
    '{name: "D28.1", is_k: 0, code_8b: 'b001_11100, code_10b_p: 'b1001_011100, code_10b_n: 'b1001_011100, flip_rd: 0},
    '{name: "D28.2", is_k: 0, code_8b: 'b010_11100, code_10b_p: 'b1010_011100, code_10b_n: 'b1010_011100, flip_rd: 0},
    '{name: "D28.3", is_k: 0, code_8b: 'b011_11100, code_10b_p: 'b0011_011100, code_10b_n: 'b1100_011100, flip_rd: 0},
    '{name: "D28.4", is_k: 0, code_8b: 'b100_11100, code_10b_p: 'b1011_011100, code_10b_n: 'b0100_011100, flip_rd: 1},
    '{name: "D28.5", is_k: 0, code_8b: 'b101_11100, code_10b_p: 'b0101_011100, code_10b_n: 'b0101_011100, flip_rd: 0},
    '{name: "D28.6", is_k: 0, code_8b: 'b110_11100, code_10b_p: 'b0110_011100, code_10b_n: 'b0110_011100, flip_rd: 0},
    '{name: "D28.7", is_k: 0, code_8b: 'b111_11100, code_10b_p: 'b0111_011100, code_10b_n: 'b1000_011100, flip_rd: 1},
    '{name: "D29.0", is_k: 0, code_8b: 'b000_11101, code_10b_p: 'b0010_011101, code_10b_n: 'b1101_100010, flip_rd: 0},
    '{name: "D29.1", is_k: 0, code_8b: 'b001_11101, code_10b_p: 'b1001_011101, code_10b_n: 'b1001_100010, flip_rd: 1},
    '{name: "D29.2", is_k: 0, code_8b: 'b010_11101, code_10b_p: 'b1010_011101, code_10b_n: 'b1010_100010, flip_rd: 1},
    '{name: "D29.3", is_k: 0, code_8b: 'b011_11101, code_10b_p: 'b1100_011101, code_10b_n: 'b0011_100010, flip_rd: 1},
    '{name: "D29.4", is_k: 0, code_8b: 'b100_11101, code_10b_p: 'b0100_011101, code_10b_n: 'b1011_100010, flip_rd: 0},
    '{name: "D29.5", is_k: 0, code_8b: 'b101_11101, code_10b_p: 'b0101_011101, code_10b_n: 'b0101_100010, flip_rd: 1},
    '{name: "D29.6", is_k: 0, code_8b: 'b110_11101, code_10b_p: 'b0110_011101, code_10b_n: 'b0110_100010, flip_rd: 1},
    '{name: "D29.7", is_k: 0, code_8b: 'b111_11101, code_10b_p: 'b1000_011101, code_10b_n: 'b0111_100010, flip_rd: 0},
    '{name: "D30.0", is_k: 0, code_8b: 'b000_11110, code_10b_p: 'b0010_011110, code_10b_n: 'b1101_100001, flip_rd: 0},
    '{name: "D30.1", is_k: 0, code_8b: 'b001_11110, code_10b_p: 'b1001_011110, code_10b_n: 'b1001_100001, flip_rd: 1},
    '{name: "D30.2", is_k: 0, code_8b: 'b010_11110, code_10b_p: 'b1010_011110, code_10b_n: 'b1010_100001, flip_rd: 1},
    '{name: "D30.3", is_k: 0, code_8b: 'b011_11110, code_10b_p: 'b1100_011110, code_10b_n: 'b0011_100001, flip_rd: 1},
    '{name: "D30.4", is_k: 0, code_8b: 'b100_11110, code_10b_p: 'b0100_011110, code_10b_n: 'b1011_100001, flip_rd: 0},
    '{name: "D30.5", is_k: 0, code_8b: 'b101_11110, code_10b_p: 'b0101_011110, code_10b_n: 'b0101_100001, flip_rd: 1},
    '{name: "D30.6", is_k: 0, code_8b: 'b110_11110, code_10b_p: 'b0110_011110, code_10b_n: 'b0110_100001, flip_rd: 1},
    '{name: "D30.7", is_k: 0, code_8b: 'b111_11110, code_10b_p: 'b1000_011110, code_10b_n: 'b0111_100001, flip_rd: 0},
    '{name: "D31.0", is_k: 0, code_8b: 'b000_11111, code_10b_p: 'b0010_110101, code_10b_n: 'b1101_001010, flip_rd: 0},
    '{name: "D31.1", is_k: 0, code_8b: 'b001_11111, code_10b_p: 'b1001_110101, code_10b_n: 'b1001_001010, flip_rd: 1},
    '{name: "D31.2", is_k: 0, code_8b: 'b010_11111, code_10b_p: 'b1010_110101, code_10b_n: 'b1010_001010, flip_rd: 1},
    '{name: "D31.3", is_k: 0, code_8b: 'b011_11111, code_10b_p: 'b1100_110101, code_10b_n: 'b0011_001010, flip_rd: 1},
    '{name: "D31.4", is_k: 0, code_8b: 'b100_11111, code_10b_p: 'b0100_110101, code_10b_n: 'b1011_001010, flip_rd: 0},
    '{name: "D31.5", is_k: 0, code_8b: 'b101_11111, code_10b_p: 'b0101_110101, code_10b_n: 'b0101_001010, flip_rd: 1},
    '{name: "D31.6", is_k: 0, code_8b: 'b110_11111, code_10b_p: 'b0110_110101, code_10b_n: 'b0110_001010, flip_rd: 1},
    '{name: "D31.7", is_k: 0, code_8b: 'b111_11111, code_10b_p: 'b1000_110101, code_10b_n: 'b0111_001010, flip_rd: 0},

    '{name: "K28.0", is_k: 1, code_8b: 'b000_11100, code_10b_p: 'b0010_111100, code_10b_n: 'b1101_000011, flip_rd: 0},
    '{name: "K28.1", is_k: 1, code_8b: 'b001_11100, code_10b_p: 'b1001_111100, code_10b_n: 'b0110_000011, flip_rd: 1},
    '{name: "K28.2", is_k: 1, code_8b: 'b010_11100, code_10b_p: 'b1010_111100, code_10b_n: 'b0101_000011, flip_rd: 1},
    '{name: "K28.3", is_k: 1, code_8b: 'b011_11100, code_10b_p: 'b1100_111100, code_10b_n: 'b0011_000011, flip_rd: 1},
    '{name: "K28.4", is_k: 1, code_8b: 'b100_11100, code_10b_p: 'b0100_111100, code_10b_n: 'b1011_000011, flip_rd: 0},
    '{name: "K28.5", is_k: 1, code_8b: 'b101_11100, code_10b_p: 'b0101_111100, code_10b_n: 'b1010_000011, flip_rd: 1},
    '{name: "K28.6", is_k: 1, code_8b: 'b110_11100, code_10b_p: 'b0110_111100, code_10b_n: 'b1001_000011, flip_rd: 1},
    '{name: "K28.7", is_k: 1, code_8b: 'b111_11100, code_10b_p: 'b0001_111100, code_10b_n: 'b1110_000011, flip_rd: 0},
    '{name: "K23.7", is_k: 1, code_8b: 'b111_10111, code_10b_p: 'b0001_010111, code_10b_n: 'b1110_101000, flip_rd: 0},
    '{name: "K27.7", is_k: 1, code_8b: 'b111_11011, code_10b_p: 'b0001_011011, code_10b_n: 'b1110_100100, flip_rd: 0},
    '{name: "K29.7", is_k: 1, code_8b: 'b111_11101, code_10b_p: 'b0001_011101, code_10b_n: 'b1110_100010, flip_rd: 0},
    '{name: "K30.7", is_k: 1, code_8b: 'b111_11110, code_10b_p: 'b0001_011110, code_10b_n: 'b1110_100001, flip_rd: 0}
  };


endpackage 