


//--------------------------------------------------------------------------
package uart_pkg;
    `timescale 1ns/1ps;

    `include "uart_base.svh";
    `include "uart_master.svh";
    `include "uart_slave.svh";

endpackage