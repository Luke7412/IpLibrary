

package axi4_pkg;

  `include "axi4_base.svh"
  `include "axi4_monitor.svh"
  `include "axi4_master.svh"
  `include "axi4_slave.svh"

endpackage