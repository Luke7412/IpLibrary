//------------------------------------------------------------------------------
// Project Name: IpLibrary
//------------------------------------------------------------------------------
// Author      : Lukas Vinkx (lvin)
// Description : 
//------------------------------------------------------------------------------


package axi4lite_pkg;

  `include "axi4lite_base.svh"
  `include "Axi4lite_Transaction.svh"
  `include "axi4lite_monitor.svh"
  `include "axi4lite_master.svh"
  `include "axi4lite_slave.svh"

endpackage