
--------------------------------------------------------------------------------
-- Info
--------------------------------------------------------------------------------
-- Hash (MD5): 0x${hash_value}
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- LIBRARIES
--------------------------------------------------------------------------------
library IEEE;
   use IEEE.STD_LOGIC_1164.ALL;


--------------------------------------------------------------------------------
-- PACKAGE HEADER
--------------------------------------------------------------------------------
package ModuleId is
   
   constant Id : std_logic_vector(127 downto 0) := X"${hash_value}";

end package;